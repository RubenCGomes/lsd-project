library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity RegInput is
	port (clk		 	: in  std_logic;
		  reset			: in  std_logic;
		  switch	 	: in  std_logic;
		  start_stop 	: in  std_logic
	);
end RegInput;

architecture Shell of RegInput is
begin

end Shell;
