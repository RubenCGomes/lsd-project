library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

entity SimpleDecounter is
	port (
	);
end SimpleDecounter;

architecture Behavioral of SimpleDecounter is
begin

end Behavioral;
